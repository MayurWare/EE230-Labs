19D070070 | Mayur Ware
*BJT Series Regulator - Analysis
*Importing the Zener Model
.SUBCKT ZENER_5.6 1 2
D1 1 2 DF
DZ 3 1 DR
VZ 2 3 4
.MODEL DF D ( IS=27.5p RS=0.620 N=1.10 CJO=78.3p VJ=1.00 M=0.330 TT=50.1n )
.MODEL DR D ( IS=5.49f RS=50 N=1.77 )
.ENDS


*Importing the SL100 and BC547
.model bc547a NPN IS=10f BF=200 ISE=10.3f IKF=50m NE=1.3
+ BR=9.5 VAF=80 IKR=12m ISC=47p NC=2 VAR=10 RB=280 RE=1 RC=40
+ tr=0.3u tf=0.5n cje=12p vje=0.48 mje=0.5 cjc=6p vjc=0.7 mjc=0.33 kf=2f
.model SL100 NPN IS=100f BF=80 ISE=10.3f IKF=50m NE=1.3
+ BR=9.5 VAF=80 IKR=12m ISC=47p NC=2 VAR=10 RB=100 RE=1 RC=10
+ tr=0.3u tf=0.5n cje=12p vje=0.48 mje=0.5 cjc=6p vjc=0.7 mjc=0.33 kf=2f

*Netlist
Rc In 1 1k
Rl Out GND 1k
X1 GND 3 ZENER_5.6
R1 Out 2 11k
R2 2 GND 14k

*Voltage Sources
Vin In GND dc 20V
 
*BJTs
Q1 In 1 Out SL100
Q2 1 2 3 bc547a

*Control Commands
.dc Vin 15 25 0.5
.control
run
set color0 = white
set color1 = black
set color2 = blue
set color3 = red
set xbrushwidth = 2
plot V(Out) V(1) V(2) V(3)
.endc
.end