RC Integrator Circuit
*Capacitor connected between In and Out
C1 In Out 0.1u 
*Resistor connected between Out and GND
R1 Out GND 10k
*Voltage Source between In and GND
Vin In GND pulse(0 5 0 0 0 10m 20m)
.tran 0.1m 100m
*Control Commands
.control
run
set color0 = white
set color1 = black
set color2 = blue
set color3 = red
set xbrushwidth = 2
plot V(In) V(Out)
.endc
.end