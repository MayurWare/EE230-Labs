19D070070 | Mayur Ware
*Common-Emitter Amplifier: Biasing Circuit
.model bc547a NPN IS=10f BF=200 ISE=10.3f IKF=50m NE=1.3
+ BR=9.5 VAF=80 IKR=12m ISC=47p NC=2 VAR=10 RB=280 RE=1 RC=40
+ tr=0.3u tf=0.5n cje=12p vje=0.48 mje=0.5 cjc=6p vjc=0.7 mjc=0.33 kf=2f
*BJT
Q1 2 3 5 bc547a
*Voltage Sources
Vin In GND 12
V1 1 2 0
V2 4 3 0
*Resistors
R1 In 4 10k
R2 4 GND 2.2k
Rc In 1 1.2k
Re 5 GND 1k
*Control Commands
.op
.control
run
print i(V2) i(V1) V(2) V(3) V(5)
.endc
.end
