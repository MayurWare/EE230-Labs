19D070070 | Mayur Ware
*Two-stage Amplifier (CE and CC): Biasing Circuit
.model bc547a NPN IS=10f BF=200 ISE=10.3f IKF=50m NE=1.3
+ BR=9.5 VAF=80 IKR=12m ISC=47p NC=2 VAR=10 RB=280 RE=1 RC=40
+ tr=0.3u tf=0.5n cje=12p vje=0.48 mje=0.5 cjc=6p vjc=0.7 mjc=0.33 kf=2f
vb2 c b2 0
ve2 e2 8 0
rc 4 3 1.2k
re 1 0 1k
r1 4 2 10k
r2 2 0 2.2k
vcc 4 0 dc 12
vb 2 b 0
vc 3 c 0
ve e 1 0 
ce 1 0 100u
c1 5 2 10u
c2 8 9 10u
re2 8 0 10k
rl 9 0 10k
vin 5 0 dc 0 ac 10m
Q1 c b e bc547a
Q2 4 b2 e2 bc547a
*Control Commands
.op
.control
run
set color0 = white
set color1 = black
set color2 = blue
set color3 = red
set xbrushwidth = 2
print V(9)
.endc
.end
