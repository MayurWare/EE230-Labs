19D070070 | Mayur Ware
*BJT Current Mirror Circuit
.model bc547a NPN IS=10f BF=100 ISE=10.3f IKF=50m NE=1.3
+ BR=9.5 VAF=200 IKR=12m ISC=47p NC=2 VAR=10 RB=280 RE=1 RC=40
+ tr=0.3u tf=0.5n cje=12p vje=0.48 mje=0.5 cjc=6p vjc=0.7 mjc=0.33 kf=2f
*BJT
Q1 2 3 GND bc547a
Q2 5 3 GND bc547a
*Voltage Sources
Vcc 1 GND 12
Vo 4 GND 1
V1 4 5 dc 0
V2 2 3 dc 0
*Resistors
R 1 2 10k
*Control Commands
.dc Vo 1 5 0.5
.control
run
set color0 = white
set color1 = black
set color2 = blue
set color3 = red
set xbrushwidth = 2
plot i(V1) 
.endc
.end