RC Integrator Circuit
*Resistor connected between In and Out
R1 In Out 10k 
*Capacitor connected between Out and GND
C1 Out GND 0.1u
*Voltage Source between In and GND
Vin In GND pulse(0 5 0 0 0 1m 2m)
.tran 0.1m 10m
*Control Commands
.control
run
set color0 = white
set color1 = black
set color2 = blue
set color3 = red
set xbrushwidth = 2
plot V(In) V(Out)
.endc
.end