19D070070 | Mayur Ware
*Two-stage Amplifier (CE and CC): Biasing Circuit
.model bc547a NPN IS=10f BF=200 ISE=10.3f IKF=50m NE=1.3
+ BR=9.5 VAF=80 IKR=12m ISC=47p NC=2 VAR=10 RB=280 RE=1 RC=40
+ tr=0.3u tf=0.5n cje=12p vje=0.48 mje=0.5 cjc=6p vjc=0.7 mjc=0.33 kf=2f
*BJT
Q1 1 2 3 bc547a
Q2 In 5 6 bc547a
*Voltage Sources
Vin In GND dc 12
V1 8 GND dc 0 ac 0.01
V2 1 5 dc 0V
V3 6 7 dc 0V
*Resistors
R1 In 2 10k
R2 2 GND 2.2k
Rc In 1 1.2k
Re 3 GND 1k
Re2 7 GND 10k
Rl Out GND 10k
*Capacitors
C1 2 8 10u
C2 6 Out 10u
Ce 3 GND 100u
*Control Commands
.ac dec 10 10 10Meg
.control
run
set color0 = white
set color1 = black
set color2 = blue
set color3 = red
set xbrushwidth = 2
*print i(V2) i(V3) V(6)
plot -V(Out)*100
.endc
.end
